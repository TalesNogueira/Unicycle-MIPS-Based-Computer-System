module FPGA_Output (input wire FLAG_output, input wire [31:0] FPGA_output, output reg [7:0] decimals);
	
endmodule 